library ieee;
use ieee.std_logic_1164.all;

entity ROArch128 is
    port(input128		 	 	: in std_logic_vector(127 downto 0);
			resetComp				: in std_logic;
			chain_reset_bit 		: in std_logic; 
			boardTemp				: in std_logic_vector (6 downto 0);
			O					 	: out std_logic_vector(127 downto 0));
end entity;


architecture behav of ROArch128 is

component main is
    port(	input128		 	 	: in std_logic_vector(127 downto 0);
			resetComp				: in std_logic;
			chain_reset_bit 		: in std_logic; 
			boardTemp				: in std_logic_vector (6 downto 0);
			O					 	: out std_logic);
end component;

--signal input128 					: std_logic_vector (127 downto 0) 	:= x"ABCDEF1023456ABCD897412ABCDEF532";


begin 	
	
	GEN_ROArch:
	for I in 0 to 127 generate
		ROAX	: main port map
		(input128, resetComp, chain_reset_bit, boardTemp, O(I));
	end generate GEN_ROArch;
	
	


end architecture;