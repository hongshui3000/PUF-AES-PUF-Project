										   library ieee;
use ieee.std_logic_1164.all;

entity mux128_1 is
    port(input 			: in std_logic_vector(127 downto 0);
		 BoardSelect 	: in std_logic_vector(6 downto 0);
		 output 		: out std_logic);
--		 muxReady	  	: out std_logic);
end entity;


architecture behav of mux128_1 is
begin
	
with BoardSelect select
    output	 	<= input(0) when "0000000",
       			   input(1) when "0000001",
						input(2) when "0000010",
         		   input(3) when "0000011",
						input(4) when "0000100",
						input(5) when "0000101",
						input(6) when "0000110",
						input(7) when "0000111",
						input(8) when "0001000",
						input(9) when "0001001",
						input(10) when "0001010",
						input(11) when "0001011",
						input(12) when "0001100",
         		   input(13) when "0001101",
						input(14) when "0001110",
						input(15) when "0001111",
						input(16) when "0010000",
						input(17) when "0010001",
						input(18) when "0010010",
						input(19) when "0010011",
						input(20) when "0010100",
						input(21) when "0010101",
						input(22) when "0010110",
         		   input(23) when "0010111",
						input(24) when "0011000",
						input(25) when "0011001",
						input(26) when "0011010",
						input(27) when "0011011",
						input(28) when "0011100",
						input(29) when "0011101",
						input(30) when "0011110",
						input(31) when "0011111",
						input(32) when "0100000",
         		   input(33) when "0100001",
						input(34) when "0100010",
						input(35) when "0100011",
						input(36) when "0100100",
						input(37) when "0100101",
						input(38) when "0100110",
						input(39) when "0100111",
						input(40) when "0101000",
						input(41) when "0101001",
						input(42) when "0101010",						
						input(43) when "0101011",
						input(44) when "0101100",
						input(45) when "0101101",	
						input(46) when "0101110",
						input(47) when "0101111",
						input(48) when "0110000",
						input(49) when "0110001",
						input(50) when "0110010",
						input(51) when "0110011",							
						input(52) when "0110100",						
						input(53) when "0110101",							
						input(54) when "0110110",						
						input(55) when "0110111",							
						input(56) when "0111000",						
						input(57) when "0111001",							
						input(58) when "0111010",						
						input(59) when "0111011",							
						input(60) when "0111100",						
						input(61) when "0111101",							
						input(62) when "0111110",						
						input(63) when "0111111",							
						input(64) when "1000000",						
						input(65) when "1000001",							
						input(66) when "1000010",						
						input(67) when "1000011",							
						input(68) when "1000100",						
						input(69) when "1000101",							
						input(70) when "1000110",						
						input(71) when "1000111",							
						input(72) when "1001000",						
						input(73) when "1001001",							
						input(74) when "1001010",						
						input(75) when "1001011",							
						input(76) when "1001100",						
						input(77) when "1001101",							
						input(78) when "1001110",						
						input(79) when "1001111",							
						input(80) when "1010000",						
						input(81) when "1010001",							
						input(82) when "1010010",						
						input(83) when "1010011",							
						input(84) when "1010100",						
						input(85) when "1010101",							
						input(86) when "1010110",						
						input(87) when "1010111",							
						input(88) when "1011000",						
						input(89) when "1011001",							
						input(90) when "1011010",
						input(91) when "1011011",							
						input(92) when "1011100",						
						input(93) when "1011101",							
						input(94) when "1011110",						
						input(95) when "1011111",							
						input(96) when "1100000",						
						input(97) when "1100001",							
						input(98) when "1100010",						
						input(99) when "1100011",							
						input(100) when "1100100",						
						input(101) when "1100101",							
						input(102) when "1100110",						
						input(103) when "1100111",							
						input(104) when "1101000",						
						input(105) when "1101001",							
						input(106) when "1101010",						
						input(107) when "1101011",							
						input(108) when "1101100",						
						input(109) when "1101101",							
						input(110) when "1101110",
						input(111) when "1101111",							
						input(112) when "1110000",						
						input(113) when "1110001",							
						input(114) when "1110010",						
						input(115) when "1110011",							
						input(116) when "1110100",						
						input(117) when "1110101",							
						input(118) when "1110110",						
						input(119) when "1110111",							
						input(120) when "1111000",						
						input(121) when "1111001",							
						input(122) when "1111010",						
						input(123) when "1111011",							
						input(124) when "1111100",						
						input(125) when "1111101",							
						input(126) when "1111110",						
						input(127) when "1111111",							
					
         		   '0'  when others;	
--with BoardSelect select
--	muxReady 	<= '1' when "0000000",
--       			   '1' when "0000001",
--						'1' when "0000010",
--         		   '1' when "0000011",
--						'1' when "0000100",
--						'1' when "0000101",
--						'1' when "0000110",
--						'1' when "0000111",
--						'1' when "0001000",
--						'1' when "0001001",
--						'1' when "0001010",
--						'1' when "0001011",
--						'1' when "0001100",
--         		   '1' when "0001101",
--						'1' when "0001110",
--						'1' when "0001111",
--						'1' when "0010000",
--						'1' when "0010001",
--						'1' when "0010010",
--						'1' when "0010011",
--						'1' when "0010100",
--						'1' when "0010101",
--						'1' when "0010110",
--         		   '1' when "0010111",
--						'1' when "0011000",
--						'1' when "0011001",
--						'1' when "0011010",
--						'1' when "0011011",
--						'1' when "0011100",
--						'1' when "0011101",
--						'1' when "0011110",
--						'1' when "0011111",
--						'1' when "0100000",
--         		   '1' when "0100001",
--						'1' when "0100010",
--						'1' when "0100011",
--						'1' when "0100100",
--						'1' when "0100101",
--						'1' when "0100110",
--						'1' when "0100111",
--						'1' when "0101000",
--						'1' when "0101001",
--						'1' when "0101010",						
--						'1' when "0101011",
--						'1' when "0101100",
--						'1' when "0101101",	
--						'1' when "0101110",
--						'1' when "0101111",
--						'1' when "0110000",
--						'1' when "0110001",
--						'1' when "0110010",
--						'1' when "0110011",							
--						'1' when "0110100",						
--						'1' when "0110101",							
--						'1' when "0110110",						
--						'1' when "0110111",							
--						'1' when "0111000",						
--						'1' when "0111001",							
--						'1' when "0111010",						
--						'1' when "0111011",							
--						'1' when "0111100",						
--						'1' when "0111101",							
--						'1' when "0111110",						
--						'1' when "0111111",							
--						'1' when "1000000",						
--						'1' when "1000001",							
--						'1' when "1000010",						
--						'1' when "1000011",							
--						'1' when "1000100",						
--						'1' when "1000101",							
--						'1' when "1000110",						
--						'1' when "1000111",							
--						'1' when "1001000",						
--						'1' when "1001001",							
--						'1' when "1001010",						
--						'1' when "1001011",							
--						'1' when "1001100",						
--						'1' when "1001101",							
--						'1' when "1001110",						
--						'1' when "1001111",							
--						'1' when "1010000",						
--						'1' when "1010001",							
--						'1' when "1010010",						
--						'1' when "1010011",							
--						'1' when "1010100",						
--						'1' when "1010101",							
--						'1' when "1010110",						
--						'1' when "1010111",							
--						'1' when "1011000",						
--						'1' when "1011001",							
--						'1' when "1011010",
--						'1' when "1011011",							
--						'1' when "1011100",						
--						'1' when "1011101",							
--						'1' when "1011110",						
--						'1' when "1011111",							
--						'1' when "1100000",						
--						'1' when "1100001",							
--						'1' when "1100010",						
--						'1' when "1100011",							
--						'1' when "1100100",						
--						'1' when "1100101",							
--						'1' when "1100110",						
--						'1' when "1100111",							
--						'1' when "1101000",						
--						'1' when "1101001",							
--						'1' when "1101010",						
--						'1' when "1101011",							
--						'1' when "1101100",						
--						'1' when "1101101",							
--						'1' when "1101110",
--						'1' when "1101111",							
--						'1' when "1110000",						
--						'1' when "1110001",							
--						'1' when "1110010",						
--						'1' when "1110011",							
--						'1' when "1110100",						
--						'1' when "1110101",							
--						'1' when "1110110",						
--						'1' when "1110111",							
--						'1' when "1111000",						
--						'1' when "1111001",							
--						'1' when "1111010",						
--						'1' when "1111011",							
--						'1' when "1111100",						
--						'1' when "1111101",							
--						'1' when "1111110",						
--						'1' when "1111111",
--						
--         		   '0'  when others;	
--				   			   
end architecture;